//////////////////////////////////////////////////////////////////////////////////
// Exercise #3 - Active IoT Devices Monitor
// Student Name:
// Date: 
//
//  Description: In this exercise, you need to design a counter of active IoT devices, where 
//  if the rst=1, the counter should be set to zero. If event=0, the value
//  should stay constant. If on-off=1, the counter should count up every
//  clock cycle, otherwise it should count down.
//  Wrap-around values are allowed.
//
//  inputs:
//           clk, rst, change, on_off
//
//  outputs:
//           counter_out[7:0]
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

module monitor (
    //Todo: add ports 
	input clk,
	input rst,
	input change,
	input on_off,
	output counter_out[7:0]

    );
                    
    //Todo: add registers and wires, if needed
//variables
wire c
wire d
always @(posedge clk) begin
	c +=1
	d -= 1
end

    //Todo: add user logic
	AND2(clk,on_off)
        assign counter_out = (rst==0) ? 0:
	assign counter_out = (on_off==1) ? c
	assign counter_out = (on_off == 0) ? d

endmodule
